class in_sequence extends  uvm_sequence;
		// component utils
	`uvm_object_utils(in_sequence)
	// class constructor function
	function void new ();
		
	endfunction : new	
	
endclass : in_sequence