class in_driver extends  uvm_component;
	// component utils
	`uvm_componnet_utils(fifo_config)
	// class constructor function
	function void new ();
		
	endfunction : new	
	
endclass : in_driver