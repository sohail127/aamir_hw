class in_agent extends  uvm_agent;
	// component utils
	`uvm_component_utils(in_agent)
	// class constructor function
	function void new ();
		
	endfunction : new

endclass : in_agent