package spi_test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  // import spi_pkg::*;
  // import spi_tb_pkg::*;


  // tests here
  `include "spi_base_test.sv"
endpackage : spi_test_pkg
