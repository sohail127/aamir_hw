`timescale 1ns/1ps
//********************************************************************************
// Title       : PUF ro
// Project     : ASIC Implementation of PUF
//********************************************************************************
// File        : puf_ro.v
// Author      : sohail (Email: sohail@imse-cnm.csic.es)
// Company     : IMSE-CNM (http://www.imse-cnm.csic.es)
// Created     : Tue Apr 12 16:33:24 2022
// Standard    : Verilog 2012
//********************************************************************************
// Copyright (c) 2022 IMSE-CNME ()
//********************************************************************************
// Description:
//********************************************************************************

module tb_puf_ro ();

//********************************************************************************
// ** Parameters declaration
//********************************************************************************
	parameter N_STAGE=5;

//********************************************************************************
// ** Inputs are reg
//********************************************************************************
	reg i_en ;
//********************************************************************************
// ** outputs are wire
//********************************************************************************
	wire o_ro;
//********************************************************************************
// ** DUT instantiation
//********************************************************************************

puf_ro #(.N_STAGE(N_STAGE)) DUT (
	.i_en(i_en), //input  i_en,
	.o_ro(o_ro)  //output o_ro
);

//********************************************************************************
// ** initzation task
//********************************************************************************
task init_sys();
	i_en = 1'b1;
endtask // init_sys

//********************************************************************************
// procedural block
//********************************************************************************
initial begin
	$display("**********************************************");
	$display("********Start Simulation**********************");
	$display("**********************************************");
	init_sys();
	#200;
	$display("**********************************************");	
	$display("********Simulation Done***********************");
	$display("**********************************************");
	$stop;
end

endmodule // tb_puf_ro