class spi_seq_pkg extends  /* base class*/;
	
endclass : spi_seq_pkg