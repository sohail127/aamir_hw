package spi_tb_pkg;
    // import uvm package and macros
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  import spi_pkg::*;

  `include "spi_env.sv"

endpackage: spi_tb_pkg