module spi();
endmodule 
