class fifo_config extends  uvm_object;
	// component utils
	`uvm_object_utils(fifo_config)
	// class constructor function
	function void new ();
		
	endfunction : new	
	
endclass : fifo_config