module sp_ram (
  input clk,    // Clock
  input clk_en, // Clock Enable
  input rst_n,  // Asynchronous reset active low
  
);

// read logic here

endmodule : sp_ram