module puf_soc_ro_decoder #(parameter MUX_LENGTH = 16) (
	input 															clk 			 ,
	input                               rst_n      ,
	input                               i_dcod_en  ,
	input      [$clog2(MUX_LENGTH)-1:0] i_sel_mux_0,
	input      [$clog2(MUX_LENGTH)-1:0] i_sel_mux_1,
	output reg [        MUX_LENGTH-1:0] o_puf_en    
);
	always@(posedge clk or negedge rst_n) begin
		if (!rst_n) begin
			o_puf_en <= {MUX_LENGTH{1'b0}};
		end else begin
			if (i_dcod_en) begin
				case (i_sel_mux_0)
					4'd0 : begin
						case (i_sel_mux_1)
							4'd1    : o_puf_en <= 16'b0000_0000_0000_0011;
							4'd2    : o_puf_en <= 16'b0000_0000_0000_0101;
							4'd3    : o_puf_en <= 16'b0000_0000_0000_1001;
							4'd4    : o_puf_en <= 16'b0000_0000_0001_0001;
							4'd5    : o_puf_en <= 16'b0000_0000_0010_0001;
							4'd6    : o_puf_en <= 16'b0000_0000_0100_0001;
							4'd7    : o_puf_en <= 16'b0000_0000_1000_0001;
							4'd8    : o_puf_en <= 16'b0000_0001_0000_0001;
							4'd9    : o_puf_en <= 16'b0000_0010_0000_0001;
							4'd10   : o_puf_en <= 16'b0000_0100_0000_0001;
							4'd11   : o_puf_en <= 16'b0000_1000_0000_0001;
							4'd12   : o_puf_en <= 16'b0001_0000_0000_0001;
							4'd13   : o_puf_en <= 16'b0010_0000_0000_0001;
							4'd14   : o_puf_en <= 16'b0100_0000_0000_0001;
							4'd15   : o_puf_en <= 16'b1000_0000_0000_0001;
							default : o_puf_en <= 16'b0000_0000_0000_0001;
						endcase
					end
					4'd1 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_0000_0011;
							4'd2    : o_puf_en <= 16'b0000_0000_0000_0110;
							4'd3    : o_puf_en <= 16'b0000_0000_0000_1010;
							4'd4    : o_puf_en <= 16'b0000_0000_0001_0010;
							4'd5    : o_puf_en <= 16'b0000_0000_0010_0010;
							4'd6    : o_puf_en <= 16'b0000_0000_0100_0010;
							4'd7    : o_puf_en <= 16'b0000_0000_1000_0010;
							4'd8    : o_puf_en <= 16'b0000_0001_0000_0010;
							4'd9    : o_puf_en <= 16'b0000_0010_0000_0010;
							4'd10   : o_puf_en <= 16'b0000_0100_0000_0010;
							4'd11   : o_puf_en <= 16'b0000_1000_0000_0010;
							4'd12   : o_puf_en <= 16'b0001_0000_0000_0010;
							4'd13   : o_puf_en <= 16'b0010_0000_0000_0010;
							4'd14   : o_puf_en <= 16'b0100_0000_0000_0010;
							4'd15   : o_puf_en <= 16'b1000_0000_0000_0010;
							default : o_puf_en <= 16'b0000_0000_0000_0010;
						endcase
					end
					4'd2 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_0000_0101;
							4'd1    : o_puf_en <= 16'b0000_0000_0000_0110;
							4'd3    : o_puf_en <= 16'b0000_0000_0000_1100;
							4'd4    : o_puf_en <= 16'b0000_0000_0001_0100;
							4'd5    : o_puf_en <= 16'b0000_0000_0010_0100;
							4'd6    : o_puf_en <= 16'b0000_0000_0100_0100;
							4'd7    : o_puf_en <= 16'b0000_0000_1000_0100;
							4'd8    : o_puf_en <= 16'b0000_0001_0000_0100;
							4'd9    : o_puf_en <= 16'b0000_0010_0000_0100;
							4'd10   : o_puf_en <= 16'b0000_0100_0000_0100;
							4'd11   : o_puf_en <= 16'b0000_1000_0000_0100;
							4'd12   : o_puf_en <= 16'b0001_0000_0000_0100;
							4'd13   : o_puf_en <= 16'b0010_0000_0000_0100;
							4'd14   : o_puf_en <= 16'b0100_0000_0000_0100;
							4'd15   : o_puf_en <= 16'b1000_0000_0000_0100;
							default : o_puf_en <= 16'b0000_0000_0000_0100;
						endcase
					end
					4'd3 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_0000_1001;
							4'd1    : o_puf_en <= 16'b0000_0000_0000_1010;
							4'd2    : o_puf_en <= 16'b0000_0000_0000_1100;
							4'd4    : o_puf_en <= 16'b0000_0000_0001_1000;
							4'd5    : o_puf_en <= 16'b0000_0000_0010_1000;
							4'd6    : o_puf_en <= 16'b0000_0000_0100_1000;
							4'd7    : o_puf_en <= 16'b0000_0000_1000_1000;
							4'd8    : o_puf_en <= 16'b0000_0001_0000_1000;
							4'd9    : o_puf_en <= 16'b0000_0010_0000_1000;
							4'd10   : o_puf_en <= 16'b0000_0100_0000_1000;
							4'd11   : o_puf_en <= 16'b0000_1000_0000_1000;
							4'd12   : o_puf_en <= 16'b0001_0000_0000_1000;
							4'd13   : o_puf_en <= 16'b0010_0000_0000_1000;
							4'd14   : o_puf_en <= 16'b0100_0000_0000_1000;
							4'd15   : o_puf_en <= 16'b1000_0000_0000_1000;
							default : o_puf_en <= 16'b0000_0000_0000_1000;
						endcase
					end
					4'd4 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_0001_0001;
							4'd1    : o_puf_en <= 16'b0000_0000_0001_0010;
							4'd2    : o_puf_en <= 16'b0000_0000_0001_0100;
							4'd3    : o_puf_en <= 16'b0000_0000_0001_1000;
							4'd5    : o_puf_en <= 16'b0000_0000_0011_0000;
							4'd6    : o_puf_en <= 16'b0000_0000_0101_0000;
							4'd7    : o_puf_en <= 16'b0000_0000_1001_0000;
							4'd8    : o_puf_en <= 16'b0000_0001_0001_0000;
							4'd9    : o_puf_en <= 16'b0000_0010_0001_0000;
							4'd10   : o_puf_en <= 16'b0000_0100_0001_0000;
							4'd11   : o_puf_en <= 16'b0000_1000_0001_0000;
							4'd12   : o_puf_en <= 16'b0001_0000_0001_0000;
							4'd13   : o_puf_en <= 16'b0010_0000_0001_0000;
							4'd14   : o_puf_en <= 16'b0100_0000_0001_0000;
							4'd15   : o_puf_en <= 16'b1000_0000_0001_0000;
							default : o_puf_en <= 16'b0000_0000_0001_0000;
						endcase
					end
					4'd5 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_0010_0001;
							4'd1    : o_puf_en <= 16'b0000_0000_0010_0010;
							4'd2    : o_puf_en <= 16'b0000_0000_0010_0100;
							4'd3    : o_puf_en <= 16'b0000_0000_0010_1000;
							4'd4    : o_puf_en <= 16'b0000_0000_0011_0000;
							4'd6    : o_puf_en <= 16'b0000_0000_0110_0000;
							4'd7    : o_puf_en <= 16'b0000_0000_1010_0000;
							4'd8    : o_puf_en <= 16'b0000_0001_0010_0000;
							4'd9    : o_puf_en <= 16'b0000_0010_0010_0000;
							4'd10   : o_puf_en <= 16'b0000_0100_0010_0000;
							4'd11   : o_puf_en <= 16'b0000_1000_0010_0000;
							4'd12   : o_puf_en <= 16'b0001_0000_0010_0000;
							4'd13   : o_puf_en <= 16'b0010_0000_0010_0000;
							4'd14   : o_puf_en <= 16'b0100_0000_0010_0000;
							4'd15   : o_puf_en <= 16'b1000_0000_0010_0000;
							default : o_puf_en <= 16'b0000_0000_0010_0000;
						endcase
					end
					4'd6 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_0100_0001;
							4'd1    : o_puf_en <= 16'b0000_0000_0100_0010;
							4'd2    : o_puf_en <= 16'b0000_0000_0100_0100;
							4'd3    : o_puf_en <= 16'b0000_0000_0100_1000;
							4'd4    : o_puf_en <= 16'b0000_0000_0101_0000;
							4'd5    : o_puf_en <= 16'b0000_0000_0110_0000;
							4'd7    : o_puf_en <= 16'b0000_0000_1100_0000;
							4'd8    : o_puf_en <= 16'b0000_0001_0100_0000;
							4'd9    : o_puf_en <= 16'b0000_0010_0100_0000;
							4'd10   : o_puf_en <= 16'b0000_0100_0100_0000;
							4'd11   : o_puf_en <= 16'b0000_1000_0100_0000;
							4'd12   : o_puf_en <= 16'b0001_0000_0100_0000;
							4'd13   : o_puf_en <= 16'b0010_0000_0100_0000;
							4'd14   : o_puf_en <= 16'b0100_0000_0100_0000;
							4'd15   : o_puf_en <= 16'b1000_0000_0100_0000;
							default : o_puf_en <= 16'b0000_0000_0100_0000;
						endcase
					end
					4'd7 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0000_1000_0001;
							4'd1    : o_puf_en <= 16'b0000_0000_1000_0010;
							4'd2    : o_puf_en <= 16'b0000_0000_1000_0100;
							4'd3    : o_puf_en <= 16'b0000_0000_1000_1000;
							4'd4    : o_puf_en <= 16'b0000_0000_1001_0000;
							4'd5    : o_puf_en <= 16'b0000_0000_1010_0000;
							4'd6    : o_puf_en <= 16'b0000_0000_1100_0000;
							4'd8    : o_puf_en <= 16'b0000_0001_1000_0000;
							4'd9    : o_puf_en <= 16'b0000_0010_1000_0000;
							4'd10   : o_puf_en <= 16'b0000_0100_1000_0000;
							4'd11   : o_puf_en <= 16'b0000_1000_1000_0000;
							4'd12   : o_puf_en <= 16'b0001_0000_1000_0000;
							4'd13   : o_puf_en <= 16'b0010_0000_1000_0000;
							4'd14   : o_puf_en <= 16'b0100_0000_1000_0000;
							4'd15   : o_puf_en <= 16'b1000_0000_1000_0000;
							default : o_puf_en <= 16'b0000_0000_1000_0000;
						endcase
					end
					4'd8 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0001_0000_0001;
							4'd1    : o_puf_en <= 16'b0000_0001_0000_0010;
							4'd2    : o_puf_en <= 16'b0000_0001_0000_0100;
							4'd3    : o_puf_en <= 16'b0000_0001_0000_1000;
							4'd4    : o_puf_en <= 16'b0000_0001_0001_0000;
							4'd5    : o_puf_en <= 16'b0000_0001_0010_0000;
							4'd6    : o_puf_en <= 16'b0000_0001_0100_0000;
							4'd7    : o_puf_en <= 16'b0000_0001_1000_0000;
							4'd9    : o_puf_en <= 16'b0000_0011_0000_0000;
							4'd10   : o_puf_en <= 16'b0000_0101_0000_0000;
							4'd11   : o_puf_en <= 16'b0000_1001_0000_0000;
							4'd12   : o_puf_en <= 16'b0001_0001_0000_0000;
							4'd13   : o_puf_en <= 16'b0010_0001_0000_0000;
							4'd14   : o_puf_en <= 16'b0100_0001_0000_0000;
							4'd15   : o_puf_en <= 16'b1000_0001_0000_0000;
							default : o_puf_en <= 16'b0000_0001_0000_0000;
						endcase
					end
					4'd9 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0010_0000_0001;
							4'd1    : o_puf_en <= 16'b0000_0010_0000_0010;
							4'd2    : o_puf_en <= 16'b0000_0010_0000_0100;
							4'd3    : o_puf_en <= 16'b0000_0010_0000_1000;
							4'd4    : o_puf_en <= 16'b0000_0010_0001_0000;
							4'd5    : o_puf_en <= 16'b0000_0010_0010_0000;
							4'd6    : o_puf_en <= 16'b0000_0010_0100_0000;
							4'd7    : o_puf_en <= 16'b0000_0010_1000_0000;
							4'd8    : o_puf_en <= 16'b0000_0011_0000_0000;
							4'd10   : o_puf_en <= 16'b0000_0110_0000_0000;
							4'd11   : o_puf_en <= 16'b0000_1010_0000_0000;
							4'd12   : o_puf_en <= 16'b0001_0010_0000_0000;
							4'd13   : o_puf_en <= 16'b0010_0010_0000_0000;
							4'd14   : o_puf_en <= 16'b0100_0010_0000_0000;
							4'd15   : o_puf_en <= 16'b1000_0010_0000_0000;
							default : o_puf_en <= 16'b0000_0010_0000_0000;
						endcase
					end
					4'd10 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_0100_0000_0001;
							4'd1    : o_puf_en <= 16'b0000_0100_0000_0010;
							4'd2    : o_puf_en <= 16'b0000_0100_0000_0100;
							4'd3    : o_puf_en <= 16'b0000_0100_0000_1000;
							4'd4    : o_puf_en <= 16'b0000_0100_0001_0000;
							4'd5    : o_puf_en <= 16'b0000_0100_0010_0000;
							4'd6    : o_puf_en <= 16'b0000_0100_0100_0000;
							4'd7    : o_puf_en <= 16'b0000_0100_1000_0000;
							4'd8    : o_puf_en <= 16'b0000_0101_0000_0000;
							4'd9    : o_puf_en <= 16'b0000_0110_0000_0000;
							4'd11   : o_puf_en <= 16'b0000_1100_0000_0000;
							4'd12   : o_puf_en <= 16'b0001_0100_0000_0000;
							4'd13   : o_puf_en <= 16'b0010_0100_0000_0000;
							4'd14   : o_puf_en <= 16'b0100_0100_0000_0000;
							4'd15   : o_puf_en <= 16'b1000_0100_0000_0000;
							default : o_puf_en <= 16'b0000_0100_0000_0000;
						endcase
					end
					4'd11 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0000_1000_0000_0001;
							4'd1    : o_puf_en <= 16'b0000_1000_0000_0010;
							4'd2    : o_puf_en <= 16'b0000_1000_0000_0100;
							4'd3    : o_puf_en <= 16'b0000_1000_0000_1000;
							4'd4    : o_puf_en <= 16'b0000_1000_0001_0000;
							4'd5    : o_puf_en <= 16'b0000_1000_0010_0000;
							4'd6    : o_puf_en <= 16'b0000_1000_0100_0000;
							4'd7    : o_puf_en <= 16'b0000_1000_1000_0000;
							4'd8    : o_puf_en <= 16'b0000_1001_0000_0000;
							4'd9    : o_puf_en <= 16'b0000_1010_0000_0000;
							4'd10   : o_puf_en <= 16'b0000_1100_0000_0000;
							4'd12   : o_puf_en <= 16'b0001_1000_0000_0000;
							4'd13   : o_puf_en <= 16'b0010_1000_0000_0000;
							4'd14   : o_puf_en <= 16'b0100_1000_0000_0000;
							4'd15   : o_puf_en <= 16'b1000_1000_0000_0000;
							default : o_puf_en <= 16'b0000_1000_0000_0000;
						endcase
					end
					4'd12 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0001_0000_0000_0001;
							4'd1    : o_puf_en <= 16'b0001_0000_0000_0010;
							4'd2    : o_puf_en <= 16'b0001_0000_0000_0100;
							4'd3    : o_puf_en <= 16'b0001_0000_0000_1000;
							4'd4    : o_puf_en <= 16'b0001_0000_0001_0000;
							4'd5    : o_puf_en <= 16'b0001_0000_0010_0000;
							4'd6    : o_puf_en <= 16'b0001_0000_0100_0000;
							4'd7    : o_puf_en <= 16'b0001_0000_1000_0000;
							4'd8    : o_puf_en <= 16'b0001_0001_0000_0000;
							4'd9    : o_puf_en <= 16'b0001_0010_0000_0000;
							4'd10   : o_puf_en <= 16'b0001_0100_0000_0000;
							4'd11   : o_puf_en <= 16'b0001_1000_0000_0000;
							4'd13   : o_puf_en <= 16'b0011_0000_0000_0000;
							4'd14   : o_puf_en <= 16'b0101_0000_0000_0000;
							4'd15   : o_puf_en <= 16'b1001_0000_0000_0000;
							default : o_puf_en <= 16'b0001_0000_0000_0000;
						endcase
					end
					4'd13 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0010_0000_0000_0001;
							4'd1    : o_puf_en <= 16'b0010_0000_0000_0010;
							4'd2    : o_puf_en <= 16'b0010_0000_0000_0100;
							4'd3    : o_puf_en <= 16'b0010_0000_0000_1000;
							4'd4    : o_puf_en <= 16'b0010_0000_0001_0000;
							4'd5    : o_puf_en <= 16'b0010_0000_0010_0000;
							4'd6    : o_puf_en <= 16'b0010_0000_0100_0000;
							4'd7    : o_puf_en <= 16'b0010_0000_1000_0000;
							4'd8    : o_puf_en <= 16'b0010_0001_0000_0000;
							4'd9    : o_puf_en <= 16'b0010_0010_0000_0000;
							4'd10   : o_puf_en <= 16'b0010_0100_0000_0000;
							4'd11   : o_puf_en <= 16'b0010_1000_0000_0000;
							4'd12   : o_puf_en <= 16'b0011_0000_0000_0000;
							4'd14   : o_puf_en <= 16'b0110_0000_0000_0000;
							4'd15   : o_puf_en <= 16'b1010_0000_0000_0000;
							default : o_puf_en <= 16'b0010_0000_0000_0000;
						endcase
					end
					4'd14 : begin
						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b0100_0000_0000_0001;
							4'd1    : o_puf_en <= 16'b0100_0000_0000_0010;
							4'd2    : o_puf_en <= 16'b0100_0000_0000_0100;
							4'd3    : o_puf_en <= 16'b0100_0000_0000_1000;
							4'd4    : o_puf_en <= 16'b0100_0000_0001_0000;
							4'd5    : o_puf_en <= 16'b0100_0000_0010_0000;
							4'd6    : o_puf_en <= 16'b0100_0000_0100_0000;
							4'd7    : o_puf_en <= 16'b0100_0000_1000_0000;
							4'd8    : o_puf_en <= 16'b0100_0001_0000_0000;
							4'd9    : o_puf_en <= 16'b0100_0010_0000_0000;
							4'd10   : o_puf_en <= 16'b0100_0100_0000_0000;
							4'd11   : o_puf_en <= 16'b0100_1000_0000_0000;
							4'd12   : o_puf_en <= 16'b0101_0000_0000_0000;
							4'd13   : o_puf_en <= 16'b0110_0000_0000_0000;
							4'd15   : o_puf_en <= 16'b1100_0000_0000_0000;
							default : o_puf_en <= 16'b0100_0000_0000_0000;
						endcase
					end
					4'd15 : begin

						case (i_sel_mux_1)
							4'd0    : o_puf_en <= 16'b1000_0000_0000_0001;
							4'd1    : o_puf_en <= 16'b1000_0000_0000_0010;
							4'd2    : o_puf_en <= 16'b1000_0000_0000_0100;
							4'd3    : o_puf_en <= 16'b1000_0000_0000_1000;
							4'd4    : o_puf_en <= 16'b1000_0000_0001_0000;
							4'd5    : o_puf_en <= 16'b1000_0000_0010_0000;
							4'd6    : o_puf_en <= 16'b1000_0000_0100_0000;
							4'd7    : o_puf_en <= 16'b1000_0000_1000_0000;
							4'd8    : o_puf_en <= 16'b1000_0001_0000_0000;
							4'd9    : o_puf_en <= 16'b1000_0010_0000_0000;
							4'd10   : o_puf_en <= 16'b1000_0100_0000_0000;
							4'd11   : o_puf_en <= 16'b1000_1000_0000_0000;
							4'd12   : o_puf_en <= 16'b1001_0000_0000_0000;
							4'd13   : o_puf_en <= 16'b1010_0000_0000_0000;
							4'd14   : o_puf_en <= 16'b1100_0000_0000_0000;
							default : o_puf_en <= 16'b1000_0000_0000_0000;
						endcase
					end
					default : o_puf_en <= 16'b0000_0000_0000_0000;
				endcase
			end else begin
				o_puf_en <= o_puf_en;
				// o_puf_en = 16'b0000_0000_0000_0000;
			end
		end
	end

endmodule // 