module shift_register #(parameter BUS_WIDTH=32) (
	input                  clk       , // clock
	input                  rst_n     , // active low reset
	input                  i_ld_data , // 1: to load data
	input                  i_sht_lr  , // shift_lr : 1 for right shift, 0: for left shift
	input  [BUS_WIDTH-1:0] i_reg_data, // register data
	output                 o_busy    , // 1: when shifiting
	output                 o_shift   , // serial output
	output                 o_valid     // 1: when output is valid
);

	// register declaration
	reg [BUS_WIDTH-1:0] reg_data   ;
	reg                 reg_o_shift;
	reg                 reg_o_busy ;
	reg                 reg_o_valid;
	reg                 reg_o_shift;
	// load and shift logic here
	always@*(posedge clk) begin
		if (!rst_n) begin
			reg_data    <= {BUS_WIDTH{1'b0}};
			reg_o_busy  <= 1'b0;
			reg_o_valid <= 1'b0;
			reg_o_shift <= 1'b0;
		end
		else	begin
			if (i_ld_data) begin
				o_reg_data <= i_reg_data;
			end
			else	begin
				if (i_sht_lr) begin // 1: for righr shift
					reg_o_shift <= reg_data[0];
					reg_data    <= {1'b0,reg_data[BUS_WIDTH-1:1]}; // right shift
					reg_o_busy  <= 1'b1;
					reg_o_valid <= 1'b1;
				end
				else	begin
					reg_o_shift <= reg_data[BUS_WIDTH-1];
					reg_data    <= {reg_data[BUS_WIDTH-1:1],1'b0}; // right left
					reg_o_busy  <= 1'b1;
					reg_o_valid <= 1'b1;
				end
			end
		end
	end

	assign o_busy  = reg_o_busy  ;
	assign o_valid = reg_o_valid ;
	assign o_shift = reg_o_shift ;

endmodule