	interface puf_tx_if (input clk); 
	logic i_tx_ready ;
	logic o_tx_data ;
	logic o_tx_valid;
endinterface : puf_tx_if