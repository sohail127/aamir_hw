`timescale 1ns/1ps
//********************************************************************************
// Title       : PUF ro
// Project     : ASIC Implementation of PUF
//********************************************************************************
// File        : puf_ro.v
// Author      : sohail (Email: sohail@imse-cnm.csic.es)
// Company     : IMSE-CNM (http://www.imse-cnm.csic.es)
// Created     : Tue Apr 12 16:33:24 2022
// Standard    : Verilog 2012
//********************************************************************************
// Copyright (c) 2022 IMSE-CNME ()
//********************************************************************************
// Description:
//********************************************************************************

module tb_puf_soc_ro_bank ();

//********************************************************************************
// ** Parameters declaration
//********************************************************************************
	parameter PUF_LENGTH   = 16;
	parameter NO_PUF_STAGE = 24;
//********************************************************************************
// ** Inputs are reg
//********************************************************************************
	reg [PUF_LENGTH-1:0] i_puf_en;
//********************************************************************************
// ** outputs are wire
//********************************************************************************
	wire [PUF_LENGTH-1:0] o_puf_ro;
//********************************************************************************
// ** DUT instantiation
//********************************************************************************

	puf_soc_ro_bank #(
		.PUF_LENGTH  (PUF_LENGTH  ),
		.NO_PUF_STAGE(NO_PUF_STAGE)
	) DUT (
		.i_puf_en(i_puf_en), // input  [PUF_LENGTH-1:0] i_puf_en, // i_puf_en
		.o_puf_ro(o_puf_ro)  // output [PUF_LENGTH-1:0] o_puf_ro
	);

//********************************************************************************
// ** initzation task
//********************************************************************************
	task init_sys();
		i_puf_en = {$bits(i_puf_en){1'b0}};
		#10
		i_puf_en = 16'b0000_0000_1000_0001;
	endtask// init_sys

//********************************************************************************
// procedural block
//********************************************************************************
	initial begin
		$display("**********************************************");
		$display("********Start Simulation**********************");
		$display("**********************************************");
		init_sys();
		#200;
		$display("**********************************************");
		$display("********Simulation Done***********************");
		$display("**********************************************");
		$stop;
	end

endmodule // tb_puf_soc_ro_bank