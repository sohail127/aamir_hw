class in_seq_item extends  uvm_object;
	// component utils
	`uvm_object_utils(in_seq_item)
	// class constructor function
	function void new ();
		
	endfunction : new	
	
endclass : in_seq_item