class in_monitor extends  uvm_monitor;
	// component utils
	`uvm_component_utils(in_monitor)
	// class constructor function
	function void new ();
		
	endfunction : new		
	
endclass : in_monitor