
class out_monitor extends  uvm_agent;
	// component utils
	`uvm_component_utils(out_monitor)
	// class constructor function
	function void new ();
		
	endfunction : new

endclass : out_monitor