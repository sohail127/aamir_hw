class fifo_base_test extends  uvm_test;
	// component utils
	`uvm_component_utils(fifo_base_test)
	// class constructor function
	function void new ();
		
	endfunction : new	
		
endclass : fifo_base_test