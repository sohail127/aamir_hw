class fifo_coverage extends  uvm_subscriber;
	// component utils
	`uvm_component_utils(fifo_config)
	// class constructor function
	function void new ();
		
	endfunction : new	
		
endclass : fifo_coverage