class in_sqr extends  uvm_sequencer;
		// component utils
	`uvm_component_utils(in_sqr)
	// class constructor function
	function void new ();
		
	endfunction : new
endclass : in_sqr