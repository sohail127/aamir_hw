class host_item;
	// data members
	int challenge_q [$] ;
	int rspns ; 
	rand int challenge ;
endclass : host_item