class out_agent extends  uvm_agent;
	
	// component utils
	`uvm_component_utils(out_agent)
	// class constructor function
	function void new ();
		
	endfunction : new

endclass : out_agent